// This file is nedded for EDAplayground
`include "generator.sv"
`include "drivers.sv"
`include "monitors.sv"
`include "agents.sv"
`include "scoreboard.sv"
`include "env.sv"
`include "test.sv"
`include "tb.sv"

