// This file is needed for EDAplayground
`include "decoders.sv"
`include "synchronizer.sv"
`include "wr_ctrl.sv"
`include "rd_ctrl.sv"
`include "fifo_mem.sv"
`include "g_fifo_if.sv"
`include "g_fifo.sv"

